`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Tianjin University
// Engineer: xlxlqqq
// 
// Create Date: 2021/06/16 08:37:32
// Design Name: 
// Module Name: Syn_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Syn_top(
    input clk,
    input rst_n,
    input button_REG,
    
    output reg [4:0] cs_pin_1
    );


 
endmodule
